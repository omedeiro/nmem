* Template netlist for nmem cell read simulation
* Generated from LTspice 24.1.4 for Windows.
I1 0 N001 PWL file=ENABPWL
I2 0 N003 PWL file=CHANPWL
R1 N001 N002 1n
R2 N003 out 1n
R3 out 0 50
R4 out 0 1G
X§HL N002 N004 out 0 tempL N005 N007 hTron_behav chan_width=250n, chan_length=2.2u, heater_resistance=150
X§HR N004 0 out 0 tempR N006 N008 hTron_behav chan_width=350n, chan_length=4u, heater_resistance=300
R§irhr N008 0 1
R§ichr N006 0 1
R§irhl N007 0 1
R§ichl N005 0 1
.tran {start_time} {stop_time} {start_save} {time_step}
.options reltol 1e-6
.lib hTron_behavioral.lib
.backanno
.end
