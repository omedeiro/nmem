I1 0 N001 400µ
I2 0 out PWL(0 0 100u 300u 200u 0 300u -300u 400u 0)
R1 out 0 50
R§ic N003 0 1
R§ir N004 0 1
X§hTron N002 0 out 0 temp N003 N004 hTron_behav
R2 N001 N002 1m
R3 out 0 1G
.tran 0 400u 0 1n
.options reltol 1e-6
.lib hTron_behavioral.lib
.backanno
.end
