* hTron IV Sweep Circuit Template
* Single hTron device characterization

* Current sources
I1 0 heater_in {I_heater}
I2 0 out PWL(0 0 100u {I_bias} 200u 0 300u {-I_bias} 400u 0)

* hTron device using behavioral model
X_hTron heater_in 0 out 0 temp Meas_Isw Meas_Ihs hTron_behav chan_width=100n, chan_length=4u, heater_resistance=300
* Load resistor
R1 out 0 50

* Additional measurement resistors
R§ic Meas_Isw 0 1
R§ir Meas_Ihs 0 1

* Parameters - only bias currents are variable
.param I_bias=300u I_heater=500u

* Analysis
.tran 0 85u 0 1n
.options reltol 1e-6

* Include behavioral model
.lib hTron_behavioral.lib

.end
